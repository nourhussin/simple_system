package SYS_PKG;
    typedef logic [7:0] dataframe_t;
endpackage